-- Cabeçalho ----
-- Cawan da Silveira Soares --
-- Gabriel Casali --

Library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity full_adder is
port(
x, y, c_in : in std_logic;
s, c_out : out std_logic
);
end full_adder;

architecture arq_full_adder of full_adder is

signal tempS, tempC, tempC2 : std_logic;

component half_adder
port(
a, b : in std_logic;
sum, carry: out std_logic
);
end component;

begin

Half1: half_adder
port map(a => x, b => y, sum => tempS, carry=> tempC);

Half2: half_adder
port map(a => tempS, b => c_in, sum => s, carry=>tempC2);

c_out <= tempC or tempC2;

end arq_full_adder;