-- Cawan Soares e Gabriel Casali
Library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity decodificador is
    port(
        x : in std_logic_vector(5 downto 0);
        display7_2 : out std_logic_vector(6 downto 0);
        display7_1 : out std_logic_vector(6 downto 0);
        display7_0 : out std_logic_vector(6 downto 0)
    );
end decodificador;

architecture estrutural of decodificador is
begin

	with x select  
--Unidade
 display7_0 <=
 --Positivos
	"1000000" when "000000"|"001010"|"010100"|"011110",
	"1111001" when "000001"|"001011"|"010101"|"011111",
	"0100100" when "000010"|"001100"|"010110",
	"0110000" when "000011"|"001101"|"010111",
	"0011001" when "000100"|"001110"|"011000",
	"0010010" when "000101"|"001111"|"011001",
	"0000010" when "000110"|"010000"|"011010",
	"1011000" when "000111"|"010001"|"011011",
	"0000000" when "001000"|"010010"|"011100",
	"0010000" when "001001"|"010011"|"011101",
--Negativos
	"1000000" when "110110"|"101100"|"100010", 
	"1111001" when "111111"|"110101"|"101011"|"100001", 
	"0100100" when "111110"|"110100"|"101010"|"100000", 
	"0110000" when "111101"|"110011"|"101001", 
	"0011001" when "111100"|"110010"|"101000", 
	"0010010" when "111011"|"110001"|"100111",
	"0000010" when "111010"|"110000"|"100110", 
	"1011000" when "111001"|"101111"|"100101", 
	"0000000" when "111000"|"101110"|"100100", 
	"0010000" when "110111"|"101101"|"100011",  
	"0000110" when others;
	
	with x select
--Dezenas
	display7_1 <=
--Positivos
	"1000000" when "000000"|"000001"|"000010"|"000011"|"000100"|"000101"|"000110"|"000111"|"001000"|"001001",
	"1111001" when "001010"|"001011"|"001100"|"001101"|"001110"|"001111"|"010000"|"010001"|"010010"|"010011",
	"0100100" when "010100"|"010101"|"010110"|"010111"|"011000"|"011001"|"011010"|"011011"|"011100"|"011101",
	"0110000" when "011110"|"011111",	
--Negativos
	"1000000" when "111111"|"111110"|"111101"|"111100"|"111011"|"111010"|"111001"|"111000"|"110111",
	"1111001" when "110110"|"110101"|"110100"|"110011"|"110010"|"110001"|"110000"|"101111"|"101110"|"101101",
	"0100100" when "101100"|"101011"|"101010"|"101001"|"101000"|"100111"|"100110"|"100101"|"100100"|"100011",
	"0110000" when "100010"|"100001"|"100000",
	"0000110" when others;
	
-- Sinal
	display7_2 <=
   "0111111" when x(5) = '1'
   else "1111111";
	



end estrutural;